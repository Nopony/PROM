* C:\Users\strad\Documents\University Stuff\PROM\lightbulb.asc
XU1 0 N004 N006 NC_01 P001 NC_02 N001 N002 NE555
V1 N002 0 5
R1 0 N001 500
D1 N001 N003 1N4148
D2 N003 N001 1N4148
C1 0 P001 100µF
Q1 12vPwm N005 0 0 2N2222
R2 N005 N006 500
R3 N003 N004 5K
C2 0 N004 100µF
.model D D
.lib C:\Users\strad\Documents\LTspiceXVII\lib\cmp\standard.dio
.model NPN NPN
.model PNP PNP
.lib C:\Users\strad\Documents\LTspiceXVII\lib\cmp\standard.bjt
.tran 20mS
.lib NE555.sub
.backanno
.end